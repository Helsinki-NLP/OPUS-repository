Presenterad av statsminister Göran Persson för den svenska riksdagen, 22 mars 1996
Fru talman, ärade ledamöter av Sveriges riksdag!
Att minska arbetslösheten är den främsta och allt annat överskuggande uppgiften för min regering.
Målet är att Sverige år 2000 skall ha halverat den öppna arbetslösheten till 4 procent.
Fundamenten för ett gott samhälle undergrävs av dagens höga arbetslöshet.
Såväl samhällsekonomi som moral och vilja försvagas.
Ytterst handlar kampen för sysselsättning om att hålla samman Sverige.
Regeringens politik mot arbetslösheten skall bygga på fyra hörnstenar:
Den första hörnstenen är stabila och uthålliga finanser.
Goda statsfinanser är grunden för alla politiska ambitioner.
Saneringen av de offentliga finanserna skall fortsätta.
Målet är att 1997 begränsa underskottet till mindre än tre procent av BNP och att Sverige år 1998 skall ha de offentliga finanserna i balans.
En ny budgetprocess med en starkare budgetuppföljning och nominella utgiftstak skapar goda förutsättningar att påbörja den nödvändiga minskningen av den offentliga skuldbördan.
Prisökningarna har pressats ned till under två procent.Inflationen skall bibehållas på en låg nivå.
Därmed skapas utrymme för fortsatta räntenedgångar.
Regeringen kan under inga omständigheter acceptera att välfärdssamhället återigen undermineras av stora underskott och en skenande statsskuld.
Den andra hörnstenen är goda villkor för företag och företagande.
Sverige är ett bra land för företagsamhet.
Här finns en flexibel ekonomi, ett konstruktivt samarbetsklimat och en kunnig och välutbildad arbetskraft.
Regeringen kommer att ytterligare förbättra företagandets villkor.
Antalet nya arbeten i små och medelstora företag har ökat kraftigt.
Det är en sund utveckling som skall stärkas genom kompetensutveckling, innovationsstöd, kapitalförsörjning och företagsstöd.
Regeringens samlade politik skall ge förbättrade möjligheter till nystartande, utveckling och expansion.
Näringspolitikens lokala och regionala roll skall framhävas.
Därigenom kan den regionala utvecklingen stärkas, EU:s strukturfonder utnyttjas bättre och näringslivet främjas.
