Lika lön för lika arbete är en grundläggande strävan.
Kvinnor och män skall ha samma möjligheter att försörja sig själva och kombinera ett utvecklande yrkesliv med ett aktivt föräldraskap.
Invandrarnas särskilda kompetens skall tas bättre till vara.
Därmed stärks Sveriges möjligheter i den ökande internationaliseringen.
Inom Europeiska unionen sluter nu allt fler länder upp bakom tanken att utarbeta gemensamma ambitioner för kampen mot arbetslöshet.
Det är en framgång.
För att intensifiera detta arbete är det av stor vikt att ett särskilt kapitel om sysselsättning skrivs in i EU:s fördrag.
Uthålliga statsfinanser, goda villkor för företagande, ett livslångt lärande och ett kontrakt för samverkan är de fyra hörnstenarna.
På denna grund bjuder regeringen in de politiska partierna, arbetsmarknadens parter och hela svenska folket att gemensamt betvinga arbetslösheten.
Endast så kan vi förverkliga våra bästa drömmars Sverige.
Globaliseringen och internationaliseringen har dramatiskt förändrat politikens möjligheter och människors liv.
Trygghet är inte längre bara en nationell angelägenhet.
För att lösa de stora och långsiktiga frågorna om fred, demokrati, trygghet och miljö krävs ett ökat internationellt samarbete.
Därför koncentreras politiken till fyra områden.
1.
EU-samarbetet skall bättre tas tillvara.
Sveriges medlemskap i Europeiska unionen bygger på en lång tradition av internationellt engagemang, solidaritet och samarbete.
Regeringen kommer aktivt att utnyttja de möjligheter som Sveriges medlemskap ger att skapa välfärd och gemensam säkerhet i vår del av världen.
EU-frågorna skall ges en ökad tyngd i den inrikespolitiska processen.
Den regeringskonferens om EU:s framtid som inleds om några dagar bör bana väg för EU:s utvidgning.
Därtill skall Sverige aktivt driva frågorna om minskad arbetslöshet, ökad öppenhet och god miljö.
2.
Fred, demokrati och social rättvisa skall säkras i hela världen.
Sveriges engagemang och ansvar stannar inte vid Europas gränser.
Förenta nationerna utgör det viktigaste redskapet för internationell fred och säkerhet, och för att hantera de globala hoten mot människans överlevnad.
Därför engagerar sig regeringen med kraft i FN:s akuta svårigheter och i behovet av reformer.
Sveriges kandidatur till FN:s säkerhetsråd är ett uttryck för vårt orubbliga stöd för ett effektivt internationellt samarbete.
Vi vill föra kampen vidare för social rättvisa, mänskliga rättigheter och en fortsatt nedrustning i världen.
En värld i djup obalans, ekonomiskt och socialt, blir aldrig säker.
Därför fullföljer regeringen traditionen av ett aktivt engagemang för folken i Mellanöstern, Afrika, Asien och Latinamerika.
Sveriges militära alliansfrihet, syftande till att vårt land skall kunna vara neutralt i händelse av krig i vårt närområde, består.
Alliansfriheten kombineras med ett aktivt ansvarstagande för säkerheten också i vår omvärld.
Svensk frivillig personal utför en viktig och riskfylld uppgift i Bosnien.
Genom vårt deltagande i fredsstyrkan IFOR ger Sverige ett konkret bidrag till de internationella ansträngningarna att bistå parterna i det sargade landet att uppnå en varaktig fred.
De nya demokratierna är bräckliga och utsatta för svåra påfrestningar.
De behöver vårt stöd i arbetet med att åter bygga upp sina samhällen och sina ekonomier.
Vi stärker Sverige genom att hjälpa andra.
Östersjökonferensen i Visby i maj blir ett viktigt startskott för en bred offensiv för utveckling och förnyelse runt Östersjön.
Östersjön skall åter göras till ett hav som förenar, utvecklar och berikar människor.
Därigenom kan en trygg grundval för demokrati och fred skapas.
3.
Miljön skall bli en tydlig och långsiktig prioritering.
Hotet mot miljön är ett hot mot livet självt.
Regeringens ambition är att Sverige skall vara en pådrivande internationell kraft och ett föregångsland i strävan att skapa ett hållbart samhälle.
De ekologiska kraven kan leda till nästa stora språng i tillväxten.
Det krävs aktiva medborgare, men också en tydlig politik, för att främja ett ökat kretsloppstänkande.
Ett nytt energisystem skall utvecklas.
Avvecklingen av kärnkraften bör inledas under mandatperioden och därefter fortsätta i jämn takt.
Den skall ske på ett sådant sätt att den elintensiva industrins konkurrensläge inte äventyras.
På grundval av 1991 års energiöverenskommelse, Energikommissionens betänkande och remissvaren på detta inbjuds samtliga riksdagspartier till överläggningar om energipolitiken.
4.
Trygghet och ansvar skall prägla samhället.
Den svenska välfärden skall omfatta alla.
Den generella välfärden är effektiv och oöverträffad i sin förmåga att skapa rättvisa och trygghet för var och en.
Den möjliggör för människan att fullt ut använda sin vilja och sin kapacitet.
Socialförsäkringarna och bidragssystemen skall ge trygghet i en föränderlig vardag.Bidrag och försäkringar skall anpassas till det förhållande att byten av yrken, liksom byten mellan arbete, studier och egenföretagande, har blivit vanligare.
Fusk och överutnyttjande av systemen kan aldrig tolereras och skall bekämpas.
Välfärd förutsätter en rättvis fördelning.
I hela världen ser vi att orättvisor och ofärd leder till ökad kriminalitet.
Brottsligheten hotar människors trygghet och även demokratin.
Vi kan aldrig tolerera ett samhälle där rädslan breder ut sig.
Kulturen och medierna skall bidra till att klyftor kan överbryggas och till att respekten och förståelsen mellan människor kan öka.
Mångfald och mångsidighet är nödvändigt för demokratin.
Kulturarvet måste vårdas, liksom de värden som det mångkulturella Sverige skapar.
En radio och TV i allmänhetens tjänst garanterar ett programutbud som når alla.
Arbetslösheten, segregationen och rasismen är de mest oroande problemen i dagens samhälle.
Om vi inte lyckas befästa idén om alla människors lika värde riskerar samhället att brytas sönder av inre motsättningar.
Därför måste hela Sverige mobiliseras för att medverka till en ökad integration.
Det är av särskild vikt att kampen mot arbetslösheten bland invandrare ges förtur.
Arbetet för ett jämställt samhälle fortsätter.
Ett jämställdhetsperspektiv skall genomsyra alla delar av regeringens politik.
En hög kvalitet i den kommunala verksamheten är grunden för den svenska välfärden, och avgörande för jämställdheten och för att motverka segregation.
Även i fortsättningen kommer den kommunala verksamheten i vård, omsorg och skola att prioriteras framför statliga bidrag och transfereringar.
För att utbudet av kommunala tjänster skall fördelas jämnt har ett nytt system för utjämning av kostnader och inkomster mellan kommunerna införts.
Det skall noga följas upp och utvärderas.
Den uppgörelse som har slutits mellan staten, Landstingsförbundet och Kommunförbundet skapar goda förutsättningar för kommunernas verksamhet och för samhällsekonomin.
Kommunerna får stabila spelregler.
Kommunala uppsägningar och skattehöjningar motverkas.
Därigenom förbättras möjligheten att bekämpa arbetslösheten.
Sverige är ett rikt land.
Vi har en god miljö, en hög kunskapsnivå, en utpräglad jämlikhet och en stor öppenhet.
Dessa värden skall värnas och vidgas.
Människovärdet är alltid större än marknadsvärdet.
Regeringens mål är ett samhälle där alla människor har arbete, känner trygghet, delaktighet och ansvar, och där var och en får del av utvecklingens framsteg.
Så kan vi hålla samman Sverige.
Eders Majestäter, Eders Kungliga Högheter, herr talman, ledamöter av Sveriges riksdag!
Sveriges neutralitetspolitik är av avgörande betydelse för vårt lands fred och oberoende.
Den bidrar också till stabilitet och avspänning i vår del av världen.
Kring denna politik finns en bred folklig uppslutning.
Den kommer att fullföljas med kraft och konsekvens.
Kränkningar av svenskt territorium kommer aldrig att accepteras.
Armén kommer att reformeras och effektiviseras.
Det är regeringens föresats att söka breda lösningar i frågor som är av betydelse för vår nationella säkerhet.
Regeringen har välkomnat överenskommelsen mellan Förenta staterna och Sovjetunionen om att avskaffa de landbaserade medeldistanskärnvapnen.
Nu måste ansträngningarna inriktas på att bland annat minska de strategiska rustningarna och få till stånd ett fullständigt provstoppsavtal.
För detta verkar Sverige bland annat inom ramen för sexnationsinitiativet.
Regeringen kommer att fortsätta att arbeta aktivt för en kärnvapenfri zon i Norden och för en korridor fri från slagfältskärnvapen i Centraleuropa.
Genom att stödja u-ländernas ekonomiska och sociala utveckling vill regeringen bidra till att vända tillbakagången i de fattiga länderna och lindra skuldkrisen.
Biståndet skall vidare främja en framsynt hushållning med naturresurser och omsorg om miljön.
Regeringen kommer att verka för att en global FN-konferens om miljö och utveckling inkallas 1992.
