Systemadministratörshandbok
Det går inte att aktivera en licens med det här serienumret.
Svara inte på det här meddelandet.
