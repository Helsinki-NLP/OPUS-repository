Näringspolitikens lokala och regionala roll skall framhävas.
Därigenom kan den regionala utvecklingen stärkas, EU:s strukturfonder utnyttjas bättre och näringslivet främjas.
Kommunernas roll i arbetsmarknadspolitiken utvecklas.
Det är kommunerna som har kunskaperna om de lokala förutsättningarna och lösningarna.
Ekonomisk brottslighet skall bekämpas - både för att hävda samhällsmoralen och för att tillse att hederliga företagare inte drabbas av osund konkurrens.
Kapitalförsörjningen skall förbättras genom införandet av en sjätte AP-fond med stora möjligheter att placera sina tillgångar i små och medelstora företag.
Regeringen eftersträvar en stabilare och mer förutsägbar politik för att förbättra företagens investeringsmöjligheter och stärka den inhemska efterfrågan.
Den tredje hörnstenen är det livslånga lärandet.
Sverige skall konkurrera med hög kompetens, inte med låga löner.
Idén om det livslånga lärandet skall förverkligas.
Skolan, förskolan och skolbarnomsorgen skall integreras för att förbättra grundskolans första viktiga år.
Gymnasieskolans kvalitet skall höjas och den eftergymnasiala utbildningen byggas ut.
Ytterligare 100.000 personer skall få möjlighet till reguljär utbildning, varav 70.000 i vuxenutbildning.
De som hittills har fått minst del av samhällets utbildningsresurser skall prioriteras.
Arbetslösa skall få möjlighet att skaffa sig en gymnasieutbildning.
Den svenska högre utbildningen och forskningen skall även fortsättningsvis hålla världsklass.
Den tvärvetenskapliga och den tillämpade forskningen skall stärkas och forskningssamarbetet mellan EU-länderna utnyttjas fullt ut.
Genom att bygga ut högskolan över hela landet ges ett kraftfullt stöd för regional utveckling.
Det ger framtidshopp, det stimulerar näringslivet och det skapar nya jobb.
Den fjärde hörnstenen är ett nytt kontrakt för samverkan.
Samförstånd har varit basen för den stabilitet och framtidstro som så länge har präglat det svenska samhället.
Samarbete är nyckeln i kampen för full sysselsättning.
En minskad arbetslöshet måste kombineras med en inflation på god europeisk nivå.
Det kräver att både de fackliga organisationerna och arbetsgivarna tar ett unikt ansvar för förändringar i förhandlings- och lönebildningssystemet samt för arbetsrätten.
I sista hand har regering och riksdag ansvaret för stabiliteten på arbetsmarknaden.
