acl
acl:cleft
acl:relcl
advcl
advmod
amod
appos
aux
aux:pass
case
cc
ccomp
compound
compound:prt
conj
cop
csubj
csubj:pass
det
discourse
dislocated
expl
fixed
flat:name
iobj
list
mark
nmod
nmod:poss
nsubj
nsubj:pass
nummod
obj
obl
obl:agent
orphan
parataxis
punct
root
vocative
xcomp
